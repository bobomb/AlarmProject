//**********************************************************/
// Structured VLSI - Spring 2014
// Alarm Clock Project
// Mofidul Islam Jamal
// Graduate Student, Florida Atlantic University
// mjamal1@fau.edu
//**********************************************************/

module alarmclock(
  input wire clk, 
  input wire reset,
  input wire alarm_button, 
  input wire time_button,
  input wire[9:0] keypad_buttons
);
parameter SHOW_CURRENT = 2'h0;
parameter SHOW_ALARM = 2'h1;
parameter SHOW_KEYPAD = 2'h2;

//holds the current time signal 
wire [15:0] current_time;
//holds the alarm time value
reg [15:0] alarm_time;
//holds the time that is given by the keypad
wire [15:0] keypad_time;
//selector for display mux
reg [1:0] selector;
//7 segment inputs
wire[3:0] segment_0, segment_1, segment_2, segment_3;
//7 segment display outputs
wire[6:0] s0_disp, s1_disp, s2_disp, s3_disp;
//tells the keypad if we want to reset the shift register
wire keypad_reset_shift;
//pulse that occurs when the keypad gets a button press and shifts a value in
wire keypad_shift_pulse;
//values to hold the new time hour and minute values, in number:number format for 24 hr clock
reg[5:0] new_time_hr;
reg[5:0] new_time_min;
//signal to counting logic to read/set the new time from new_time_hr and new_time_min
reg new_time;
//signal generated by timing generator to let us know 1 second has passed
wire one_second;
//signal generated by timing generator to let us know that 1 minute has passed
wire one_minute;
//pulsed when its time to raise the alarm
wire sound_alarm;

comparator timing_comparator(clk, current_time, alarm_time, sound_alarm);
timinggenerator timing(clk, reset, one_second, one_minute);
countinglogic count(one_minute, reset, new_time, new_time_hr, new_time_min, current_time);
//note that display segement digit mapping is HH:MM in 24 hr format
// H(segment_0) H (segment_1) : M(segment_2) M(segment_3)
multiplexor display_multiplexor(current_time, alarm_time, keypad_time, selector, segment_0, segment_1, segment_2, segment_3);
//connect 7 segment display inputs and outputs
sevensegment s0(segment_0, s0_disp);
sevensegment s1(segment_1, s1_disp);
sevensegment s2(segment_2, s2_disp);
sevensegment s3(segment_3, s3_disp);

keypad keys(clk, keypad_buttons, keypad_reset_shift, keypad_time, keypad_shift_pulse);

initial begin
  selector = 2'b00;
end
initial begin
  //this is the output of the display muxes 4 digits
  $monitor($time," \n %c\t %c\t %c\t %c\n%c%c%c\t%c%c%c\t%c%c%c\t%c%c%c\n%c%c%c\t%c%c%c\t%c%c%c\t%c%c%c\n" ,
  s3_disp[0] ? "_" : " ", s2_disp[0] ? "_" : " ", s1_disp[0] ? "_" : " ", s0_disp[0] ? "_" : " ",
  
  s3_disp[5] ? "|" : " ", s3_disp[6] ? "_" : " ", s3_disp[1] ? "|" : " ", 
  s2_disp[5] ? "|" : " ", s2_disp[6] ? "_" : " ", s2_disp[1] ? "|" : " ", 
  s1_disp[5] ? "|" : " ", s1_disp[6] ? "_" : " ", s1_disp[1] ? "|" : " ", 
  s0_disp[5] ? "|" : " ", s0_disp[6] ? "_" : " ", s0_disp[1] ? "|" : " ",
   
  s3_disp[4] ? "|" : " ", s3_disp[3] ? "_" : " ", s3_disp[2] ? "|" : " ",
  s2_disp[4] ? "|" : " ", s2_disp[3] ? "_" : " ", s2_disp[2] ? "|" : " ",
  s1_disp[4] ? "|" : " ", s1_disp[3] ? "_" : " ", s1_disp[2] ? "|" : " ",
  s0_disp[4] ? "|" : " ", s0_disp[3] ? "_" : " ", s0_disp[2] ? "|" : " "
  
  );
end


endmodule