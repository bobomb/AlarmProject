//**********************************************************/
// Structured VLSI - Spring 2014
// Alarm Clock Project
// Mofidul Islam Jamal
// Graduate Student, Florida Atlantic University
// mjamal1@fau.edu
//**********************************************************/

module alarmclock(
  input wire clk, 
  input wire reset,
  input wire alarm_button, 
  input wire time_button,
  input wire[9:0] keypad_buttons
);
parameter DISP_SHOW_CURRENT = 2'h0;
parameter DISP_SHOW_ALARM = 2'h1;
parameter DISP_SHOW_KEYPAD = 2'h2;

//holds the current time signal 
wire [15:0] current_time;
//holds the alarm time value
reg [15:0] alarm_time;
//holds the time that is given by the keypad
wire [15:0] keypad_time;
//selector for display mux
reg [1:0] selector;
//7 segment inputs
wire[3:0] segment_0, segment_1, segment_2, segment_3;
//7 segment display outputs
wire[6:0] s0_disp, s1_disp, s2_disp, s3_disp;
//tells the keypad if we want to reset the shift register
wire keypad_reset_shift;
//pulse that occurs when the keypad gets a button press and shifts a value in
wire keypad_shift_pulse;
//holds values when combined with set_new_time to set the time in the counting logic
reg[15:0] new_time;
//signal to counting logic to read/set the new time from set_new_time_hr and set_new_time_min
reg set_new_time;
//signal generated by timing generator to let us know 1 second has passed
wire one_second;
//signal generated by timing generator to let us know that 1 minute has passed
wire one_minute;
//pulsed when its time to raise the alarm
wire sound_alarm;
//holds a counter for the 10 second pulse
reg[3:0] ten_second_counter;
//holds state machine state
reg[3:0] current_state; 
parameter STATE_CURRENT_TIME = 4'h0;
parameter  STATE_DISPLAY_KEYPAD = 4'h1;
parameter STATE_DISPLAY_ALARM = 4'h2;
//first hook up timing gen
timinggenerator timing(clk, reset, one_second, one_minute);
//then counting logic to keep current_time
countinglogic count(one_minute, reset, set_new_time, new_time, current_time);
//then comparator so we know to sound the alarm
comparator timing_comparator(clk, current_time, alarm_time, sound_alarm);
//note that display segement digit mapping is HH:MM in 24 hr format
// H(segment_0) H (segment_1) : M(segment_2) M(segment_3)
multiplexor display_multiplexor(current_time, alarm_time, keypad_time, selector, segment_0, segment_1, segment_2, segment_3);
//connect 7 segment display inputs and outputs
sevensegment s0(segment_0, s0_disp);
sevensegment s1(segment_1, s1_disp);
sevensegment s2(segment_2, s2_disp);
sevensegment s3(segment_3, s3_disp);
//last component is keypad
keypad keys(clk, keypad_buttons, keypad_reset_shift, keypad_time, keypad_shift_pulse);

initial begin
  selector = 2'b00;
  alarm_time = {4'h1, 4'h2, 4'h0, 4'h0}; //alarm time set for 12:00 by default
  ten_second_counter = 4'h0;
  current_state = STATE_CURRENT_TIME;
end

always@(reset, one_second, alarm_button, time_button, keypad_shift_pulse) begin
  //handle reset
  if(reset == 1) begin
    selector = 2'b00; //reset the display mux selector
    alarm_time = {4'h1, 4'h2, 4'h0, 4'h0}; //alarm time set for 12:00 by default
  end
  
  //main state machine
  case(current_state)
    STATE_CURRENT_TIME : begin
      //reset the set new time
      set_new_time = 0;
      
      selector = DISP_SHOW_CURRENT;
      //alarm button means show the alarm time
      if(alarm_button) begin
        current_state = STATE_DISPLAY_ALARM;
      end
      
      if(keypad_shift_pulse) begin
        current_state = STATE_DISPLAY_KEYPAD;
      end
    end
    STATE_DISPLAY_KEYPAD : begin
      selector = DISP_SHOW_KEYPAD;
      if(one_second) begin
        ten_second_counter = ten_second_counter + 1;
      end
      
      //check if time needs to be set
      if(time_button) begin
        new_time = keypad_time;
        set_new_time = 1;
        current_state = STATE_CURRENT_TIME;
      end
      
    end
    STATE_DISPLAY_ALARM : begin
      selector = DISP_SHOW_ALARM;
      if(!alarm_button) begin
        current_state = STATE_CURRENT_TIME;
      end
    end
  endcase
end

initial begin
  //this is the output of the display muxes 4 digits
  $monitor($time," \n %c\t %c\t %c\t %c\n%c%c%c\t%c%c%c\t%c%c%c\t%c%c%c\n%c%c%c\t%c%c%c\t%c%c%c\t%c%c%c\n" ,
  s3_disp[0] ? "_" : " ", s2_disp[0] ? "_" : " ", s1_disp[0] ? "_" : " ", s0_disp[0] ? "_" : " ",
  
  s3_disp[5] ? "|" : " ", s3_disp[6] ? "_" : " ", s3_disp[1] ? "|" : " ", 
  s2_disp[5] ? "|" : " ", s2_disp[6] ? "_" : " ", s2_disp[1] ? "|" : " ", 
  s1_disp[5] ? "|" : " ", s1_disp[6] ? "_" : " ", s1_disp[1] ? "|" : " ", 
  s0_disp[5] ? "|" : " ", s0_disp[6] ? "_" : " ", s0_disp[1] ? "|" : " ",
   
  s3_disp[4] ? "|" : " ", s3_disp[3] ? "_" : " ", s3_disp[2] ? "|" : " ",
  s2_disp[4] ? "|" : " ", s2_disp[3] ? "_" : " ", s2_disp[2] ? "|" : " ",
  s1_disp[4] ? "|" : " ", s1_disp[3] ? "_" : " ", s1_disp[2] ? "|" : " ",
  s0_disp[4] ? "|" : " ", s0_disp[3] ? "_" : " ", s0_disp[2] ? "|" : " "
  
  );
end


endmodule
